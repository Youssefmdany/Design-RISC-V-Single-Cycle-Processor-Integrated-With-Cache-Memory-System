module instr_mem (addr, inst);


input [31:0] addr;
output [31:0] inst;
reg [31:0] inst_mem [(2**16)-1:0]; 


assign inst = inst_mem[ addr[10:2] ];


initial begin
  
  
  
  
  
/* inst_mem[0]  = 32'b00000000101000000000000010010011;  // addi x1, x0, 10
inst_mem[1]  = 32'b00000001010000000000000100010011;  // addi x2, x0, 20
inst_mem[2]  = 32'b00000010100000000000000110010011;  // addi x3, x0, 40
inst_mem[3]  = 32'b00000101000000000000001000010011;  // addi x4, x0, 80
inst_mem[4]  = 32'b00001010000000000000001010010011;  // addi x5, x0, 160
inst_mem[5]  = 32'b00000000000100000010000000100011;  // sw x1, 0(x0)
inst_mem[6]  = 32'b00000000001000000010001000100011;  // sw x2, 4(x0)
inst_mem[7]  = 32'b00000000001100000010010000100011;  // sw x3, 8(x0)
inst_mem[8]  = 32'b00000000010000000010011000100011;  // sw x4, 12(x0)
inst_mem[9]  = 32'b00000000010100000010011000100011;  // sw x5, 12(x0)
inst_mem[10]  = 32'b00000000000000000010010100000011;  // lw x10, 0(x0)
inst_mem[11] = 32'b00000000010000000010010110000011;  // lw x11, 4(x0)
inst_mem[12] = 32'b00000000100000000010011000000011;  // lw x12, 8(x0)
inst_mem[13] = 32'b00000000110000000010011010000011;  // lw x13, 12(x0)
inst_mem[14] = 32'b00000000010000000010011000100011;  // sw x4, 12(x0) */ 
  
    inst_mem[0] = 32'h00500113;
    inst_mem[1] = 32'h00C00193;
    inst_mem[2] = 32'hFF718393;
    inst_mem[3] = 32'h0023E233;
    inst_mem[4] = 32'h0041F2B3;
    inst_mem[5] = 32'h004282B3;
    inst_mem[6] = 32'h02728863;
    inst_mem[7] = 32'h0041A233;
    inst_mem[8] = 32'h00020463;
    inst_mem[9] = 32'h00000293;
    inst_mem[10] = 32'h0023A233;
    inst_mem[11] = 32'h005203B3;
    inst_mem[12] = 32'h402383B3;
    inst_mem[13] = 32'h0471AA23;
    inst_mem[14] = 32'h06002103;
    inst_mem[15] = 32'h005104B3;
    inst_mem[16] = 32'h008001EF;
    inst_mem[17] = 32'h00100113;
    inst_mem[18] = 32'h00910133;
    inst_mem[19] = 32'h0221A023;
    inst_mem[20] = 32'h00210063;  
  
end

endmodule

